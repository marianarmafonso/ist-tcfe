.options savecurrents

* PHILIPS BJT'S
.MODEL BC557A PNP(IS=2.059E-14 ISE=2.971f ISC=1.339E-14 XTI=3 BF=227.3 BR=7.69 IKF=0.08719 IKR=0.07646 XTB=1.5 VAF=37.2 VAR=11.42 VJE=0.5912 VJC=0.1 RE=0.688 RC=0.6437 RB=1 RBM=1 IRB=1E-06 CJE=1.4E-11 CJC=1.113E-11 XCJC=0.6288 FC=0.7947 NF=1.003 NR=1.007 NE=1.316 NC=1.15 MJE=0.3572 MJC=0.3414 TF=7.046E-10 TR=1m2 ITF=0.1947 VTF=5.367 XTF=4.217 EG=1.11)
.MODEL BC547A NPN(IS=1.533E-14 ISE=7.932E-16 ISC=8.305E-14 XTI=3 BF=178.7 BR=8.628 IKF=0.1216 IKR=0.1121 XTB=1.5 VAF=69.7 VAR=44.7 VJE=0.4209 VJC=0.2 RE=0.6395 RC=0.6508 RB=1 RBM=1 IRB=1E-06 CJE=1.61E-11 CJC=4.388p XCJC=0.6193 FC=0.7762 NF=1.002 NR=1.004 NE=1.436 NC=1.207 MJE=0.3071 MJC=0.2793 TF=4.995E-10 TR=1m2 ITF=0.7021 VTF=3.523 XTF=139 EG=1.11)

Vcc vcc 0 12.0
Vin in 0 0 ac 1.0 sin(0 10m 1k)
Rin in in2 100

* input coupling capacitor
Ci in2 base 0.45m

* bias circuit
R1 vcc base 125.05k
R2 base 0 20k

* gain stage
Q1 coll base emit BC547A
Rc vcc coll 0.571k
Re emit 0 100

* bypass capacitor
Cb emit 0 4.465m


* output stage
Q2 0 coll emit2 BC557A
Rout emit2 vcc 100

* output coupling capacitor
Co emit2 out 1.806m

* load
RL out 0 8

.op
.end

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"


echo "********************************************"
echo  "Time analysis"
echo "********************************************"

tran 1e-5 1e-2
*plot v(coll)
*hardcopy vo1.ps vdb(coll)

echo "********************************************"
echo  "frequency analysis"
echo "********************************************"

ac dec 10 10 100MEG
*plot vdb(coll)
*plot vp(coll)
*hardcopy vo1f.ps vdb(coll)

*plot vdb(out)
*plot vp(out)
hardcopy vo2f.ps vdb(out)
echo vo2f_FIG

*calculate cutoff frequency
let limit = vecmax(vdb(out))-3
meas ac lower WHEN vdb(out) = limit RISE = 1
meas ac upper WHEN vdb(out) = limit CROSS = LAST


*input impedance in kohm
let zin1 = -v(in2)/vin#branch
let zin = abs(zin1[40])
hardcopy zin.ps abs(v(in2)/vin#branch/(-1000))
echo zin_FIG

*calculate merit 
let gain = vecmax(abs(v(out)/v(in)))
let bandwidth = upper - lower
let cost = 100/1000 + 1.8060e-3*1e6 + 125.05e3/1000 + 20e3/1000 + 0.571e3/1000 + 100/1000 + 4.465e-3*1e6 + 100/1000 + 0.45e-3*1e6 + 2*0.1
let merit = vecmax(abs(v(out)/v(in))) * (upper - lower) / lower / (100/1000 + 1.8060e-3*1e6 + 125.05e3/1000 + 20e3/1000 + 0.571e3/1000 + 100/1000 + 4.465e-3*1e6 + 100/1000 + 0.45e-3*1e6 + 2*0.1)

*print frequencies, impedancies, gain and merit

echo  "op_TAB1"
print gain lower upper bandwidth zin cost merit
echo  "op_END1"

quit
.endc 
