*Title: lab 2 simulation

.option savecurrents

.include ../mat/ngspice_t22.txt

.control

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

quit
.endc

.end
