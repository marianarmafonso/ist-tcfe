*Title: lab 1 simulation

.option savecurrents

*Netlist
Va 1 2 DC 5.13988034104
Id 0 4 DC 1.02475824097m

R1 6 1 1.00332071212k
R2 5 6 2.04460853047k
R3 6 7 3.08291730437k
R4 2 7 4.16061678649k
R5 4 7 3.04022345043k
R6 2 8 2.06711403452k
R7 3 0 1.03302701196k

*Vaux
Vaux 8 3 0V

*Ib and Vc
Hc 7 0 Vaux 8.16113797582k
Gb 4 5 (6,7) 7.0544535009m

.control

op

echo "********************************************"
echo  "Operating point"
echo "********************************************"

echo  "op_TAB"
print all
echo  "op_END"

.endc

.end
