*Title: lab 2 simulation

.option savecurrents

*Netlist

Vs 1 0 0.0 ac 1.0 sin(0 1 1k)
R1 1 2 1.00332071212k
R2 2 3 2.04460853047k
R3 2 5 3.08291730437k
R4 0 5 4.16061678649k
R5 5 6 3.04022345043k
R6 0 4 2.06711403452k
R7 7 8 1.03302701196k
C1 6 8 1.02475824097u

*Vaux
Vaux 4 7 0V

*Ib and Vd
Hd 5 8 Vaux 8.16113797582k
Gb 6 3 (2,5) 7.0544535009m

.op 

.ic v(6) = 8.671786V v(8) = 0

.end

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red

op

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 20e-3

hardcopy trans.ps v(1) v(6)
echo trans_FIG

echo "********************************************"
echo  "Frequency analysis"
echo "********************************************"

ac dec 1000 0.1 1MEG

hardcopy acm.ps vdb(1) vdb(6) db(v(6)-v(8)) ylabel 'magnitude (dB)'
echo acm_FIG

set units = degrees
hardcopy acp.ps vp(1) vp(6) ph(v(6)-v(8)) ylabel 'phase (degrees)'
echo acp_FIG

quit
.endc
