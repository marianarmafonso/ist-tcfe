*-----------------------------------------------------------------------------
*
* To use a subcircuit, the name must begin with 'X'.  For example:
* X1 1 2 3 4 5 uA741
*
* connections:   non-inverting input
*                |  inverting input
*                |  |  positive power supply
*                |  |  |  negative power supply
*                |  |  |  |  output
*                |  |  |  |  |
.subckt uA741    1  2  3  4  5
*
  c1   11 12 8.661E-12
  c2    6  7 30.00E-12
  dc    5 53 dx
  de   54  5 dx
  dlp  90 91 dx
  dln  92 90 dx
  dp    4  3 dx
  egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
  fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
  ga    6  0 11 12 188.5E-6
  gcm   0  6 10 99 5.961E-9
  iee  10  4 dc 15.16E-6
  hlim 90  0 vlim 1K
  q1   11  2 13 qx
  q2   12  1 14 qx
  r2    6  9 100.0E3
  rc1   3 11 5.305E3
  rc2   3 12 5.305E3
  re1  13 10 1.836E3
  re2  14 10 1.836E3
  ree  10 99 13.19E6
  ro1   8  5 50
  ro2   7 99 100
  rp    3  4 18.16E3
  vb    9  0 dc 0
  vc    3 53 dc 1
  ve   54  4 dc 1
  vlim  7  8 dc 0
  vlp  91  0 dc 40
  vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends



.options savecurrents

Vcc vcc 0 10.0
Vee vee 0 -10.0
Vin vin 0 0 ac 1.0 sin(0 10m 1k)

X1 in_volt inv_in vcc vee out uA741

* non-inverting input +
C1 vin in_volt 220n
R1 in_volt 0 1k

* inverting input -
R3 inv_in out 100k
R4 inv_in 0 1k

* load
R2 out vo 1k
C2 vo 0 110n

.op
.end

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=rgb:0/9/9
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0



op

print all


* time analysis *

tran 1e-5 1e-2
*plot v(vo)
*hardcopy vo1.ps v(vo)


* frequency analysis *

ac dec 1000 10 100MEG
*plot vdb(out)
*plot vp(out)

hardcopy vo1f.ps vdb(vo)
echo vo1f_FIG
hardcopy vo1p.ps vp(vo)*180/pi
echo vo1p_FIG

* Cut-off Frequency *

let Av_db = vdb(vo)-vdb(vin)
meas ac voltGainDB MAX Av_db
let threshold = voltGainDB-3

print threshold


meas ac lowfreq WHEN Av_db=threshold
meas ac Maxfreq MAX_AT Av_db
meas ac highfreq WHEN Av_db=threshold CROSS=LAST

let centerfreq = sqrt(lowfreq*highfreq)
print lowfreq highfreq Maxfreq centerfreq

* Out gain *

let out_m = vm(out)/vm(vin)
meas ac outGain MAX out_m
print outGain


* merit *

let gainDeviation = abs(voltGainDB - 40)
let freqDeviation = abs(centerfreq - 1k)
let cost = ((8.661e-12 + 30e-12)*1000000 + (100000 + 5305 + 5305 + 1836 + 1836 + 13190000 + 50 + 100 + 18160)/1000 + (2*0.1)) + 103 + (0.220*2)
let merit = 1/(cost*(gainDeviation + freqDeviation + 1e-6))
print gainDeviation freqDeviation cost merit


* impedance ohm *

*input impedance in ohm
let Zin = abs(v(vin)[20]/vin#branch[20]/(-1))
print Zin

*need a different setup to measure output impedance

echo  "op_TAB"
print lowfreq highfreq centerfreq outGain gainDeviation freqDeviation cost merit Zin
echo  "op_END"


quit
.endc 
